`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/23/2024 07:30:18 PM
// Design Name: 
// Module Name: Memory
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Memory(input clk, input MemRead, input MemWrite, 
input [2:0] fun3, input [5:0] addr, input [31:0] data_in, output reg [31:0] data_out);

 reg [7:0] mem [0:1023]; //each is 512 bytes
    
    always@(*) begin
        if(!(MemRead || MemWrite)) begin //fetching instruction
            data_out = {mem[(addr*4)+515],mem[(addr*4)+514],mem[(addr*4)+513],mem[(addr*4)+512]};
        end else begin
            if(MemRead)
                case(fun3) // reading  Data
                3'b000:data_out= {{24{mem[addr][7]}}, mem[addr]};      //LB
                3'b001:data_out={{16{mem[addr+1][7]}},mem[addr+1],mem[addr]};      //LH
                3'b010:data_out={mem[addr+3],mem[addr+2],mem[addr+1],mem[addr]};      //LW
                3'b100:data_out= {24'b0, mem[addr]};    //LBU
                3'b101:data_out={16'b0, mem[addr+1],mem[addr]};      //LHU
                default:data_out=0;
                endcase
            else data_out = 0; // dont read
        end
    end
    
    
    always@(posedge clk) begin
            if(MemWrite) begin
                case(fun3)
                        3'b000: mem[addr]<=data_in[7:0]; //SB
                        3'b001:   {mem[addr+1],mem[addr]}<=data_in[15:0]; //SH
                        3'b010:   {mem[addr+3],mem[addr+2],mem[addr+1],mem[addr]}<=data_in;   //SW
                        default: mem[addr]<=data_in[7:0]; 
                 endcase
              end
                           
           end
           
           
    initial begin 

// // # Load operations
// mem[512] = 32'b00000000000000000010111000110111; // LUI x28, 2
// mem[513] = 32'b00000000000000000010111000010111; // AUIPC x28, 2
// mem[514] = 32'b00000000000000000010000010000011; // LW x1, 0(x0)
// mem[515] = 32'b00000000000000000001000100000011; // LH x2, 4(x0)
// mem[516] = 32'b00000000000000000000000110000011; // LB x3, 0(x0)
// mem[517] = 32'b00000000000000000100001000000011; // LBU x4, 0(x0)
// mem[518] = 32'b00000000000000000101001010000011; // LHU x5, 0(x0)

// //Arithmetic operations
// mem[519] = 32'b00000000001000001000001100110011; // ADD x6, x1, x2
// mem[520] = 32'b01000000001000001000001110110011; // SUB x7, x1, x2
// mem[521] = 32'b00000000001000001100010000110011; // XOR x8, x1, x2
// mem[522] = 32'b00000000001000001110010010110011; //  OR x9, x1, x2
// mem[523] = 32'b00000000001000001111010100110011; //AND x10, x1, x2

// // # Immediate operations
// mem[524] = 32'b00000000010000001000010110010011; // ADDI x11, x1, 4
// mem[525] = 32'b00000000010000001100011000010011; // XORI x12, x1, 4
// mem[526] = 32'b00000000010000001110011010010011; //  ORI x13, x1, 4
// mem[527] = 32'b00000000010000001111011100010011; // ANDI x14, x1, 4
// mem[528] = 32'b00000000010000001010011110010011; // SLTI x15, x1, 4
// mem[529] = 32'b00000000010000001011100000010011; //SLTIU x16, x1, 4

// // Shift operations
// mem[530] = 32'b00000000001000001101100010110011; // SRL x17, x1, x2
// mem[531] = 32'b01000000001000001101100100110011; // SRA x18, x1, x2
// mem[532] = 32'b01000000000100001101100110010011; // SRAI x19, x1, 1
// mem[533] = 32'b00000000001000001001101000110011; // SLL x20, x1, x2
// mem[534] = 32'b00000000000100001001101010010011; // SLLI x21, x1, 1
// mem[535] = 32'b00000000000100001101101100010011; // SRLI x22, x1, 1

// // # Set less than operations
// mem[536] = 32'b00000000001000001010101110110011; // SLT x23, x1, x2
// mem[537] = 32'b00000000001000001011110000110011; // SLTU x24, x1, x2

// // # Store operations
// mem[538] = 32'b00000000000100000010000000100011; // SW x1, 0(x0)
// mem[539] = 32'b00000000000100000000000000100011; // SB x1, 0(x0)
// mem[540] = 32'b00000000000100000001000000100011; // SH x1, 0(x0)

// // # Branch operations
// mem[541] = 32'b00000000000000000000001001100011; // BEQ x0, x0, 4
// mem[542] = 32'b00000000000111111000111110010011; // increment x31
// mem[543] = 32'b00000000001000001001001001100011; // BNE x1, x2, 4
// mem[544] = 32'b00000000000111111000111110010011; // increment x31
// mem[545] = 32'b00000000010000011100001001100011; // BLT x3, x4, 4
// mem[546] = 32'b00000000000111111000111110010011; // increment x31
// mem[547] = 32'b00000000011000101101001001100011; // BGE x5, x6, 4
// mem[548] = 32'b00000000000111111000111110010011; // increment x31
// mem[549] = 32'b00000000100000111110001001100011; // BLTU x7, x8,4
// mem[550] = 32'b00000000000111111000111110010011; //increment  x31
// mem[551] = 32'b00000000101001001111001001100011; //BGEU x9, x10 4
// mem[552] = 32'b00000000000111111000111110010011; // increment x31

// // # Jump operations
// mem[553] = 32'b00000000010000000000111011101111; // JAL x29, 4
// mem[554] = 32'b00000000000000000000111101100111; // JALR x30, 0(x0)

// // # Fence operation,Environment call and break
// mem[555] = 32'b00001111111100000000000000001111; // FENCE
// mem[556] = 32'b00000000000100000000000001110011; // EBREAK
// mem[557] = 32'b00000000000000000000000001110011; // ECALL
















//----------------------------------------------Arithmetic------------------------------------------------
    // {mem[515],mem[514],mem[513],mem[512]} = 32'b000000000000_00000_000_00001_0000011; // lb x1, 0(x0)
    // {mem[519],mem[518],mem[517],mem[516]} = 32'b000000000001_00000_000_00010_0000011; // lb x2, 1(x0)
    // {mem[523],mem[522],mem[521],mem[520]} = 32'b000000000010_00000_000_00011_0000011; // lb x3, 2(x0)
    // {mem[527],mem[526],mem[525],mem[524]} = 32'b00000000001000001000001100110011; // ADD x6, x1, x2
    // {mem[531],mem[530],mem[529],mem[528]} = 32'b00000000001000001000001100110011; // ADD x6, x1, x2
    // {mem[535],mem[534],mem[533],mem[532]} = 32'b01000000001000001000001110110011; // SUB x7, x1, x2
    // {mem[539],mem[538],mem[537],mem[536]} = 32'b00000000001000001100010000110011; // XOR x8, x1, x2
    // {mem[543],mem[542],mem[541],mem[540]} = 32'b00000000001000001110010010110011; //  OR x9, x1, x2
    // {mem[547],mem[546],mem[545],mem[544]} = 32'b00000000001000001111010100110011; //AND x10, x1, x2
    // // {mem[551],mem[550],mem[549],mem[548]} = 32'b
    // // {mem[555],mem[554],mem[553],mem[552]} = 32'b
    // // {mem[559],mem[558],mem[557],mem[556]} = 32'b


//----------------------------------------------Immediate------------------------------------------------
    // {mem[515],mem[514],mem[513],mem[512]} = 32'b000000000000_00000_000_00001_0000011; // lb x1, 0(x0)
    // {mem[519],mem[518],mem[517],mem[516]} = 32'b00000000010000001000010110010011; // ADDI x11, x1, 4
    // {mem[523],mem[522],mem[521],mem[520]} = 32'b00000000010000001100011000010011; // XORI x12, x1, 4
    // {mem[527],mem[526],mem[525],mem[524]} = 32'b00000000010000001110011010010011; //  ORI x13, x1, 4
    // {mem[531],mem[530],mem[529],mem[528]} = 32'b00000000010000001111011100010011; // ANDI x14, x1, 4
    // {mem[535],mem[534],mem[533],mem[532]} = 32'b00000000010000001010011110010011; // SLTI x15, x1, 4
    // {mem[539],mem[538],mem[537],mem[536]} = 32'b00000000010000001011100000010011; //SLTIU x16, x1, 4
    // // {mem[543],mem[542],mem[541],mem[540]} = 
    // // {mem[547],mem[546],mem[545],mem[544]} = 
    // // {mem[551],mem[550],mem[549],mem[548]} = 32'b
    // // {mem[555],mem[554],mem[553],mem[552]} = 32'b
    // // {mem[559],mem[558],mem[557],mem[556]} = 32'b

//----------------------------------------------SHIFT------------------------------------------------


    // {mem[515],mem[514],mem[513],mem[512]} = 32'b000000000000_00000_000_00001_0000011; // lb x1, 0(x0)
    // {mem[519],mem[518],mem[517],mem[516]} = 32'b000000000001_00000_000_00010_0000011; // lb x2, 1(x0)
    // {mem[523],mem[522],mem[521],mem[520]} = 32'b00000000001000001101100010110011; // SRL x17, x1, x2
    // {mem[527],mem[526],mem[525],mem[524]} = 32'b01000000001000001101100100110011; // SRA x18, x1, x2
    // {mem[531],mem[530],mem[529],mem[528]} = 32'b01000000000100001101100110010011; // SRAI x19, x1, 1
    // {mem[535],mem[534],mem[533],mem[532]} = 32'b00000000001000001001101000110011; // SLL x20, x1, x2
    // {mem[539],mem[538],mem[537],mem[536]} = 32'b00000000000100001001101010010011; // SLLI x21, x1, 1
    // {mem[543],mem[542],mem[541],mem[540]} = 32'b00000000000100001101101100010011; // SRLI x22, x1, 1

//------------------------------------------Branching-------------------------------------------------

    // {mem[515],mem[514],mem[513],mem[512]} = 32'b000000000000_00000_000_00001_0000011; // lb x1, 0(x0)
    // {mem[519],mem[518],mem[517],mem[516]} = 32'b000000000001_00000_000_00010_0000011; // lb x2, 1(x0)
    // {mem[523],mem[522],mem[521],mem[520]} = 32'b00000000000000000000001001100011; // BEQ x0, x0, 4
    // {mem[527],mem[526],mem[525],mem[524]} = 32'b00000000000111111000111110010011; // increment x31
    // {mem[531],mem[530],mem[529],mem[528]} = 32'b00000000001000001001001001100011; // BNE x1, x2, 4
    // {mem[535],mem[534],mem[533],mem[532]} = 32'b00000000000111111000111110010011; // increment x31
    // {mem[539],mem[538],mem[537],mem[536]} = 32'b00000000001000001100001001100011; // BLT x1, x2, 4
    // {mem[543],mem[542],mem[541],mem[540]} = 32'b00000000000111111000111110010011; // increment x31
    // {mem[547],mem[546],mem[545],mem[544]} = 32'b00000000001000001101001001100011; // BGE x1, x2, 4
    // {mem[551],mem[550],mem[549],mem[548]} = 32'b00000000000111111000111110010011; // increment x31
    // {mem[555],mem[554],mem[553],mem[552]} = 32'b00000000001000001110001001100011; // BLTU x1, x2,4
    // {mem[559],mem[558],mem[557],mem[556]} = 32'b00000000000111111000111110010011; // increment x31
    // {mem[563],mem[562],mem[561],mem[560]} = 32'b00000000001000001111001001100011; // BGEU x1, x2 4
    // {mem[567],mem[566],mem[565],mem[564]} = 32'b00000000000111111000111110010011; // increment x31


//----------------------------------------Testing------------------------------------------



    {mem[515],mem[514],mem[513],mem[512]} = 32'b000000000000_00000_000_00001_0000011; // lb x1, 0(x0)
    {mem[519],mem[518],mem[517],mem[516]} =32'b00000000000000000000000001110011; // ECALL











    
//    {mem[515],mem[514],mem[513],mem[512]}=32'b000000000000_00000_010_00001_0000011; // lw x1, 0(x0)
//    {mem[519],mem[518],mem[517],mem[516]}=32'b000000000100_00000_010_00010_0000011; // lw x2, 4(x0)
//    {mem[523],mem[522],mem[521],mem[520]}=32'b000000001000_00000_010_00011_0000011; // lw x3, 8(x0)
//   {mem[527],mem[526],mem[525],mem[524]}=32'b0000000_00010_00011_000_00101_0110011; // add x5, x3, x2=25
//    {mem[531],mem[530],mem[529],mem[528]} = 32'b0000000_00101_00000_010_01100_0100011; // sw x5, 12(x0)
//    {mem[535],mem[534],mem[533],mem[532]}= 32'b000000001100_00000_010_00110_0000011; // lw x6, 12(x0)
//    {mem[539],mem[538],mem[537],mem[536]}= 32'b0000000_00001_00110_111_00111_0110011; // and x7, x6, x1
    
    end
    
    
    initial begin
//    {mem[3],mem[2],mem[1],mem[0]}=32'd11;
//    {mem[7],mem[6],mem[5],mem[4]}=32'd12;
//    {mem[11],mem[10],mem[9],mem[8]}=32'd13;
mem[0]=2;
mem[1]=3;
mem[2]=5;



// //comprehensive test
// mem[0]=8'd5;
// mem[1]=8'd0;
// mem[2]=8'd0;
// mem[3]=8'd0;

// mem[4]=8'd2;
// mem[5]=8'd0;
// mem[6]=8'd0;
// mem[7]=8'd0;

// mem[8]=8'd3;
// mem[9]=8'd0;
// mem[10]=8'd0;
// mem[11]=8'd0;

// mem[12]=8'd12;
// mem[13]=8'd13;
// mem[14]=8'd14;
// mem[15]=8'd15;
// mem[16]=8'd16;
// mem[17]=8'd17;
// mem[18]=8'd18;
// mem[19]=8'd19;
// mem[20]=8'd20;
// mem[21]=8'd21;
// mem[22]=8'd22;
// mem[23]=8'd23;
// mem[24]=8'd24;
// mem[25]=8'd25;
// mem[26]=8'd26;
// mem[27]=8'd27;
// mem[28]=8'd28;
// mem[29]=8'd29;
// mem[30]=8'd30;
// mem[31]=8'd31;
// mem[32]=8'd32;
// mem[33]=8'd33;
// mem[34]=8'd34;
// mem[35]=8'd35;
// mem[36]=8'd36;
// mem[37]=8'd37;
// mem[38]=8'd38;
// mem[39]=8'd39;
// mem[40]=8'd40;
// mem[41]=8'd41;
// mem[42]=8'd42;
// mem[43]=8'd43;
// mem[44]=8'd44;
// mem[45]=8'd45;
// mem[46]=8'd46;
// mem[47]=8'd47;
// mem[48]=8'd48;
// mem[49]=8'd49;
// mem[50]=8'd50;
// mem[51]=8'd51;
// mem[52]=8'd52;
// mem[53]=8'd53;
// mem[54]=8'd54;
// mem[55]=8'd55;
// mem[56]=8'd56;
// mem[57]=8'd57;
// mem[58]=8'd58;
// mem[59]=8'd59;
// mem[60]=8'd60;
// mem[61]=8'd61;
// mem[62]=8'd62;
// mem[63]=8'd63;

    end
   
   
endmodule
