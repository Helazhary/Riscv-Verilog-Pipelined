`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/10/2024 02:09:36 PM
// Design Name: 
// Module Name: PC
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module PC(input clk,rst, input [5:0]pc_in, output reg [5:0] pc_out);
    
    always @(posedge clk or posedge rst)begin
        if(~rst)
        pc_out = pc_in;
        else
        pc_out=0;
    end

    
    
endmodule


